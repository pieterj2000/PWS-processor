 module asdf;
 
 endmodule