// Test2.v

// Generated using ACDS version 13.0 156 at 2016.12.01.12:12:17

`timescale 1 ps / 1 ps
module Test2 (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> onchip_memory2_0:reset

	Test2_onchip_memory2_0 onchip_memory2_0 (
		.clk         (clk_clk),                        //   clk1.clk
		.address     (),                               //     s1.address
		.debugaccess (),                               //       .debugaccess
		.clken       (),                               //       .clken
		.chipselect  (),                               //       .chipselect
		.write       (),                               //       .write
		.readdata    (),                               //       .readdata
		.writedata   (),                               //       .writedata
		.byteenable  (),                               //       .byteenable
		.reset       (rst_controller_reset_out_reset)  // reset1.reset
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
